// Tick clock
`define TICK #10ns; clk = 0; #10ns; clk = 1; #1ns;